
module xor2 (
    input a,
    input b,
    output y
);
    assign y = a ^ b; // XOR 逻辑
endmodule
